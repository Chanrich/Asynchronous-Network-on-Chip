library verilog;
use verilog.vl_types.all;
entity edu_tb is
end edu_tb;
