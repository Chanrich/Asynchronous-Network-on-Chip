library verilog;
use verilog.vl_types.all;
entity edu_sv_unit is
end edu_sv_unit;
