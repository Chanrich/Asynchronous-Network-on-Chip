library verilog;
use verilog.vl_types.all;
entity arbiter_block_sv_unit is
end arbiter_block_sv_unit;
