library verilog;
use verilog.vl_types.all;
entity data_split_module_sv_unit is
end data_split_module_sv_unit;
