library verilog;
use verilog.vl_types.all;
entity computation_module_tb is
end computation_module_tb;
