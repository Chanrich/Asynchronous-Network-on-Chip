library verilog;
use verilog.vl_types.all;
entity test_bench_sv_unit is
end test_bench_sv_unit;
