library verilog;
use verilog.vl_types.all;
entity node_sv_unit is
end node_sv_unit;
