library verilog;
use verilog.vl_types.all;
entity path_comp_sv_unit is
end path_comp_sv_unit;
