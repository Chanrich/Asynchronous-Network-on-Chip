library verilog;
use verilog.vl_types.all;
entity input_process_block_tb is
end input_process_block_tb;
