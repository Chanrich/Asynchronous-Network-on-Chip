library verilog;
use verilog.vl_types.all;
entity data_splitter_tb is
end data_splitter_tb;
