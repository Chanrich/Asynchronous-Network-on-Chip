library verilog;
use verilog.vl_types.all;
entity SystemVerilogCSP_sv_unit is
end SystemVerilogCSP_sv_unit;
