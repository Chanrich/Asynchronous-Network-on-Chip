library verilog;
use verilog.vl_types.all;
entity tb_module is
end tb_module;
