library verilog;
use verilog.vl_types.all;
entity input_arbiter_block is
end input_arbiter_block;
